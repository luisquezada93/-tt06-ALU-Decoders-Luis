`default_nettype none `timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;

  // Replace tt_um_example with your module name:
  tt_um_ALU_DECODERS user_project (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(1'b1),
      .VGND(1'b0),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );
//Generate stimulus for the inputs
   initial begin
    //Default Verification
    #1; 
    #1; ui_in [7:5] = 3'b111; ui_in [4:2] = 3'b111;
    //Octal Decoder
    #1; ui_in [1:0] = 2'd0; uio_in[7] = 1'b0;
    #1; ui_in [1:0] = 2'd1;
    #1; ui_in [1:0] = 2'd2;
    #1; ui_in [1:0] = 2'd3;
    //Gray Decoder
    #1; ui_in [1:0] = 2'd0; uio_in[7] = 1'b1;
    #1; ui_in [1:0] = 2'd1;
    #1; ui_in [1:0] = 2'd2;
    #1; ui_in [1:0] = 2'd3;
    // New numbers as Input
    #1; ui_in [7:5] = 3'b101; ui_in [4:2] = 3'b011;
    //Octal Decoder
    #1; ui_in [1:0] = 2'd0; uio_in[7] = 1'b0;
    #1; ui_in [1:0] = 2'd1;
    #1; ui_in [1:0] = 2'd2;
    #1; ui_in [1:0] = 2'd3;
    //Gray Decoder
    #1; ui_in [1:0] = 2'd0; uio_in[7] = 1'b1;
    #1; ui_in [1:0] = 2'd1;
    #1; ui_in [1:0] = 2'd2;
    #1; ui_in [1:0] = 2'd3;
      
    //Parar simulación
    #100;
    $stop;
    end
endmodule
